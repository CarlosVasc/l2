*V_6(t)
.options savecurrents

.include ../doc/ngspice_3.txt

.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control


echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3 uic

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

hardcopy Sim_3.eps v(V6) 


quit
.endc

.end
